// Color macros
`define BLURPLE     { 8'd88, 8'd101, 8'd242 }
`define GREY        { 8'd44, 8'd47, 8'd51 }
`define LIGHT_GREY  { 8'd54, 8'd57, 8'd63 }
`define WHITE       { 8'd255, 8'd255, 8'd255 }

// Logo macros
`define LOGO_START_Y    0
`define LOGO_END_Y      31
`define LOGO_START_X    1
`define LOGO_END_X      117

// Server font macros
`define FONT_SERVER_YMARGIN    1
`define FONT_SERVER_HEIGHT     16

// Channel font macros
`define FONT_CHANNEL_YMARGIN   1
`define FONT_CHANNEL_HEIGHT    14

// Sidebar macros
`define SIDEBAR_SERVER_Y_OFFSET   36
`define SIDEBAR_CHANNEL_Y_OFFSET  49
`define SIDEBAR_OFFSET_X          5
`define SIDEBAR_END_X             127

